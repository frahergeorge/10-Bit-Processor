module Register
(
	input wire [9:0] D,
	input wire En,
	output wire [9:0] Q
);