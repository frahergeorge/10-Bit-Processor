module Register
(
	input wire [9:0] D,
	input wire En,
	input wire CLKb,
	output wire [9:0] Q
);